LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;
use IEEE.math_real.ALL;


ENTITY test_calculpuissance IS
END test_calculpuissance;
